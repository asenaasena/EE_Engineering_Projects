--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   08:56:59 05/05/2017
-- Design Name:   
-- Module Name:   C:/Users/user/Desktop/COURSES/EE 240/lab7/VGA_color/freq_div_tb.vhd
-- Project Name:  VGA_color
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: freq_div
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
USE ieee.numeric_std.ALL;
 
ENTITY freq_div_tb IS
END freq_div_tb;
 
ARCHITECTURE behavior OF freq_div_tb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT freq_div
    PORT(
         clock : IN  std_logic;
         reset : IN  std_logic;
         slow_clk : OUT  std_logic
        );
    END COMPONENT;
    

   --Inputs
   signal clock : std_logic := '0';
   signal reset : std_logic := '0';

 	--Outputs
   signal slow_clk : std_logic;

   -- Clock period definitions
   constant clock_period : time := 10 ns;
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: freq_div PORT MAP (
          clock => clock,
          reset => reset,
          slow_clk => slow_clk
        );

   -- Clock process definitions
   clock_process :process
   begin
		clock <= '0';
		wait for clock_period/2;
		clock <= '1';
		wait for clock_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	
        
		  
		 
      wait for clock_period*10;

      -- insert stimulus here 
        reset<='1';
		wait for 10 ns;
		 reset<='0';
		wait for 100 ns;
      wait;
   end process;

END;
